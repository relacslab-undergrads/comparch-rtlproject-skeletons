parameter [5:0] ALU_SEL_ADD = 6'b100000;
parameter [5:0] ALU_SEL_SUB = 6'b010000;
parameter [5:0] ALU_SEL_CMP = 6'b001000;
parameter [5:0] ALU_SEL_AND = 6'b000100;
parameter [5:0] ALU_SEL_OR  = 6'b000010;
parameter [5:0] ALU_SEL_XOR = 6'b000001;
